// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.


module example (
  `include "partition_ports.vh"
);


`include "cl_firesim_defines.vh" // CL Defines for cl_firesim
`include "FireSim-generated.defines.vh" // CL Defines for cl_firesim generated by firesim Makefrag

logic rst_main_n_sync;
logic rst_firesim_n_sync;
logic rst_extra1_n_sync;

//--------------------------------------------0
// Start with Tie-Off of Unused Interfaces
//---------------------------------------------
// the developer should use the next set of `include
// to properly tie-off any unused interface
// The list is put in the top of the module
// to avoid cases where developer may forget to
// remove it from the end of the file

assign irq_req = 16'b0;

//-------------------------------------------------
// Wires
//-------------------------------------------------

//-------------------------------------------------
// Reset Synchronization Outer
//-------------------------------------------------
logic pre_sync_rst_n;

always_ff @(negedge resetn or posedge clk)
   if (!resetn)
   begin
      pre_sync_rst_n  <= 0;
      rst_main_n_sync <= 0;
   end
   else
   begin
      pre_sync_rst_n  <= 1;
      rst_main_n_sync <= pre_sync_rst_n;
   end

logic pre_sync_rst_n_extra1;
always_ff @(negedge resetn or posedge clk)
   if (!resetn)
   begin
      pre_sync_rst_n_extra1  <= 0;
      rst_extra1_n_sync <= 0;
   end
   else
   begin
      pre_sync_rst_n_extra1  <= 1;
      rst_extra1_n_sync <= pre_sync_rst_n_extra1;
   end

//---------------------------

logic firesim_internal_clock;

clk_wiz_0_firesim firesim_clocking
(
    // Clock out ports
    .clk_out1(firesim_internal_clock),
    // Status and control signals
    .reset(!rst_extra1_n_sync), // input reset
    .locked(),       // output locked
   // Clock in ports
    .clk_in1(clk)      // input clk_in1, expects 125 mhz
);

//-------------------------------------------------
// Reset Synchronization Inner
//-------------------------------------------------
logic pre_sync_rst_n_firesim;
always_ff @(negedge resetn or posedge firesim_internal_clock)
   if (!resetn)
   begin
      pre_sync_rst_n_firesim  <= 0;
      rst_firesim_n_sync <= 0;
   end
   else
   begin
      pre_sync_rst_n_firesim  <= 1;
      rst_firesim_n_sync <= pre_sync_rst_n_firesim;
   end

//-------------------------------------------------
// PCIe OCL AXI-L (SH to CL) Timing Flops
//-------------------------------------------------

  // Write address                                                                                                              
  logic        sh_ocl_awvalid_q;
  logic [31:0] sh_ocl_awaddr_q;
  logic        ocl_sh_awready_q;
                                                                                                                              
  // Write data                                                                                                                
  logic        sh_ocl_wvalid_q;
  logic [31:0] sh_ocl_wdata_q;
  logic [ 3:0] sh_ocl_wstrb_q;
  logic        ocl_sh_wready_q;
                                                                                                                              
  // Write response                                                                                                            
  logic        ocl_sh_bvalid_q;
  logic [ 1:0] ocl_sh_bresp_q;
  logic        sh_ocl_bready_q;
                                                                                                                              
  // Read address                                                                                                              
  logic        sh_ocl_arvalid_q;
  logic [31:0] sh_ocl_araddr_q;
  logic        ocl_sh_arready_q;
                                                                                                                              
  // Read data/response                                                                                                        
  logic        ocl_sh_rvalid_q;
  logic [31:0] ocl_sh_rdata_q;
  logic [ 1:0] ocl_sh_rresp_q;
  logic        sh_ocl_rready_q;

// clock converter for OCL connection
axi_clock_converter_oclnew ocl_clock_convert (
  .s_axi_aclk(clk),        // input wire s_axi_aclk
  .s_axi_aresetn(rst_main_n_sync),  // input wire s_axi_aresetn

  .s_axi_awaddr(CTL_S_AXI_LITE_awaddr),    // input wire [31 : 0] s_axi_awaddr
  .s_axi_awprot(3'h0),             // input wire [2 : 0] s_axi_awprot
  .s_axi_awvalid(CTL_S_AXI_LITE_awvalid),  // input wire s_axi_awvalid
  .s_axi_awready(CTL_S_AXI_LITE_awready),  // output wire s_axi_awready
  .s_axi_wdata(CTL_S_AXI_LITE_wdata),      // input wire [31 : 0] s_axi_wdata
  .s_axi_wstrb(CTL_S_AXI_LITE_wstrb),      // input wire [3 : 0] s_axi_wstrb
  .s_axi_wvalid(CTL_S_AXI_LITE_wvalid),    // input wire s_axi_wvalid
  .s_axi_wready(CTL_S_AXI_LITE_wready),    // output wire s_axi_wready
  .s_axi_bresp(CTL_S_AXI_LITE_bresp),      // output wire [1 : 0] s_axi_bresp
  .s_axi_bvalid(CTL_S_AXI_LITE_bvalid),    // output wire s_axi_bvalid
  .s_axi_bready(CTL_S_AXI_LITE_bready),    // input wire s_axi_bready
  .s_axi_araddr(CTL_S_AXI_LITE_araddr),    // input wire [31 : 0] s_axi_araddr
  .s_axi_arprot(3'h0),             // input wire [2 : 0] s_axi_arprot
  .s_axi_arvalid(CTL_S_AXI_LITE_arvalid),  // input wire s_axi_arvalid
  .s_axi_arready(CTL_S_AXI_LITE_arready),  // output wire s_axi_arready
  .s_axi_rdata(CTL_S_AXI_LITE_rdata),      // output wire [31 : 0] s_axi_rdata
  .s_axi_rresp(CTL_S_AXI_LITE_rresp),      // output wire [1 : 0] s_axi_rresp
  .s_axi_rvalid(CTL_S_AXI_LITE_rvalid),    // output wire s_axi_rvalid
  .s_axi_rready(CTL_S_AXI_LITE_rready),    // input wire s_axi_rready

  .m_axi_aclk(firesim_internal_clock),        // input wire m_axi_aclk
  .m_axi_aresetn(rst_firesim_n_sync),  // input wire m_axi_aresetn
  .m_axi_awaddr(sh_ocl_awaddr_q),    // output wire [31 : 0] m_axi_awaddr
  .m_axi_awprot(),    // output wire [2 : 0] m_axi_awprot
  .m_axi_awvalid(sh_ocl_awvalid_q),  // output wire m_axi_awvalid
  .m_axi_awready(ocl_sh_awready_q),  // input wire m_axi_awready
  .m_axi_wdata(sh_ocl_wdata_q),      // output wire [31 : 0] m_axi_wdata
  .m_axi_wstrb(sh_ocl_wstrb_q),      // output wire [3 : 0] m_axi_wstrb
  .m_axi_wvalid(sh_ocl_wvalid_q),    // output wire m_axi_wvalid
  .m_axi_wready(ocl_sh_wready_q),    // input wire m_axi_wready
  .m_axi_bresp(ocl_sh_bresp_q),      // input wire [1 : 0] m_axi_bresp
  .m_axi_bvalid(ocl_sh_bvalid_q),    // input wire m_axi_bvalid
  .m_axi_bready(sh_ocl_bready_q),    // output wire m_axi_bready
  .m_axi_araddr(sh_ocl_araddr_q),    // output wire [31 : 0] m_axi_araddr
  .m_axi_arprot(),    // output wire [2 : 0] m_axi_arprot
  .m_axi_arvalid(sh_ocl_arvalid_q),  // output wire m_axi_arvalid
  .m_axi_arready(ocl_sh_arready_q),  // input wire m_axi_arready
  .m_axi_rdata(ocl_sh_rdata_q),      // input wire [31 : 0] m_axi_rdata
  .m_axi_rresp(ocl_sh_rresp_q),      // input wire [1 : 0] m_axi_rresp
  .m_axi_rvalid(ocl_sh_rvalid_q),    // input wire m_axi_rvalid
  .m_axi_rready(sh_ocl_rready_q)    // output wire m_axi_rready
);

//-------------------------------------------------
// PCIe DMA_PCIS to FireSim Master
//-------------------------------------------------

   logic [5:0] sh_cl_dma_pcis_awid_FIRESIM;
   logic [63:0] sh_cl_dma_pcis_awaddr_FIRESIM;
   logic [7:0] sh_cl_dma_pcis_awlen_FIRESIM;
   logic [2:0] sh_cl_dma_pcis_awsize_FIRESIM;
   logic sh_cl_dma_pcis_awvalid_FIRESIM;
   logic cl_sh_dma_pcis_awready_FIRESIM;

   logic [511:0] sh_cl_dma_pcis_wdata_FIRESIM;
   logic [63:0] sh_cl_dma_pcis_wstrb_FIRESIM;
   logic sh_cl_dma_pcis_wlast_FIRESIM;
   logic sh_cl_dma_pcis_wvalid_FIRESIM;
   logic cl_sh_dma_pcis_wready_FIRESIM;

   logic [5:0] cl_sh_dma_pcis_bid_FIRESIM_wide;
   logic [3:0] cl_sh_dma_pcis_bid_FIRESIM;
   assign cl_sh_dma_pcis_bid_FIRESIM_wide = {2'b0, cl_sh_dma_pcis_bid_FIRESIM};

   logic [1:0] cl_sh_dma_pcis_bresp_FIRESIM;
   logic cl_sh_dma_pcis_bvalid_FIRESIM;
   logic sh_cl_dma_pcis_bready_FIRESIM;

   logic [5:0] sh_cl_dma_pcis_arid_FIRESIM;
   logic [63:0] sh_cl_dma_pcis_araddr_FIRESIM;
   logic [7:0] sh_cl_dma_pcis_arlen_FIRESIM;
   logic [2:0] sh_cl_dma_pcis_arsize_FIRESIM;
   logic sh_cl_dma_pcis_arvalid_FIRESIM;
   logic cl_sh_dma_pcis_arready_FIRESIM;

   logic [5:0] cl_sh_dma_pcis_rid_FIRESIM_wide;
   logic [3:0] cl_sh_dma_pcis_rid_FIRESIM;
   assign cl_sh_dma_pcis_rid_FIRESIM_wide = {2'b0, cl_sh_dma_pcis_rid_FIRESIM};

   logic [511:0] cl_sh_dma_pcis_rdata_FIRESIM;
   logic [1:0] cl_sh_dma_pcis_rresp_FIRESIM;
   logic cl_sh_dma_pcis_rlast_FIRESIM;
   logic cl_sh_dma_pcis_rvalid_FIRESIM;
   logic sh_cl_dma_pcis_rready_FIRESIM;

   assign cl_sh_dma_wr_full = 1'b0;
   assign cl_sh_dma_rd_full = 1'b0;


wire [5 : 0] DMA_S_AXI_awid_wide;
assign DMA_S_AXI_awid_wide = {2'b0, DMA_S_AXI_awid};
wire [5 : 0] DMA_S_AXI_arid_wide;
assign DMA_S_AXI_arid_wide = {2'b0, DMA_S_AXI_arid};



axi_clock_converter_512_wide wide_pcis_clock_convert (
  .s_axi_aclk(clk),          // input wire s_axi_aclk
  .s_axi_aresetn(rst_main_n_sync),    // input wire s_axi_aresetn

  .s_axi_awid(DMA_S_AXI_awid_wide),          // input wire [5 : 0] s_axi_awid
  .s_axi_awaddr(DMA_S_AXI_awaddr),      // input wire [63 : 0] s_axi_awaddr
  .s_axi_awlen(DMA_S_AXI_awlen),        // input wire [7 : 0] s_axi_awlen
  .s_axi_awsize(DMA_S_AXI_awsize),      // input wire [2 : 0] s_axi_awsize
  .s_axi_awburst(2'b1),    // input wire [1 : 0] s_axi_awburst
  .s_axi_awlock(1'b0),      // input wire [0 : 0] s_axi_awlock
  // CACHE = xx1x indicates the transcation is modifiable and
  // that the converter should pack narrow reads into wider ones
  .s_axi_awcache(4'h2),    // input wire [3 : 0] s_axi_awcache
  .s_axi_awprot(3'b0),      // input wire [2 : 0] s_axi_awprot
  .s_axi_awregion(4'b0),  // input wire [3 : 0] s_axi_awregion
  .s_axi_awqos(4'b0),        // input wire [3 : 0] s_axi_awqos
  .s_axi_awvalid(DMA_S_AXI_awvalid),    // input wire s_axi_awvalid
  .s_axi_awready(DMA_S_AXI_awready),    // output wire s_axi_awready

  .s_axi_wdata(DMA_S_AXI_wdata),        // input wire [511 : 0] s_axi_wdata
  .s_axi_wstrb(DMA_S_AXI_wstrb),        // input wire [63 : 0] s_axi_wstrb
  .s_axi_wlast(DMA_S_AXI_wlast),        // input wire s_axi_wlast
  .s_axi_wvalid(DMA_S_AXI_wvalid),      // input wire s_axi_wvalid
  .s_axi_wready(DMA_S_AXI_wready),      // output wire s_axi_wready

  .s_axi_bid(DMA_S_AXI_bid),            // output wire [5 : 0] s_axi_bid
  .s_axi_bresp(DMA_S_AXI_bresp),        // output wire [1 : 0] s_axi_bresp
  .s_axi_bvalid(DMA_S_AXI_bvalid),      // output wire s_axi_bvalid
  .s_axi_bready(DMA_S_AXI_bready),      // input wire s_axi_bready

  .s_axi_arid(DMA_S_AXI_arid_wide),          // input wire [5 : 0] s_axi_arid
  .s_axi_araddr(DMA_S_AXI_araddr),      // input wire [63 : 0] s_axi_araddr
  .s_axi_arlen(DMA_S_AXI_arlen),        // input wire [7 : 0] s_axi_arlen
  .s_axi_arsize(DMA_S_AXI_arsize),      // input wire [2 : 0] s_axi_arsize
  .s_axi_arburst(2'b1),    // input wire [1 : 0] s_axi_arburst
  .s_axi_arlock(1'b0),      // input wire [0 : 0] s_axi_arlock
  // CACHE = xx1x indicates the transcation is modifiable and
  // that the converter should pack narrow reads into wider ones
  .s_axi_arcache(4'h2),    // input wire [3 : 0] s_axi_arcache
  .s_axi_arprot(3'b0),      // input wire [2 : 0] s_axi_arprot
  .s_axi_arregion(4'b0),  // input wire [3 : 0] s_axi_arregion
  .s_axi_arqos(4'b0),        // input wire [3 : 0] s_axi_arqos
  .s_axi_arvalid(DMA_S_AXI_arvalid),    // input wire s_axi_arvalid
  .s_axi_arready(DMA_S_AXI_arready),    // output wire s_axi_arready

  .s_axi_rid(DMA_S_AXI_rid),            // output wire [5 : 0] s_axi_rid
  .s_axi_rdata(DMA_S_AXI_rdata),        // output wire [511 : 0] s_axi_rdata
  .s_axi_rresp(DMA_S_AXI_rresp),        // output wire [1 : 0] s_axi_rresp
  .s_axi_rlast(DMA_S_AXI_rlast),        // output wire s_axi_rlast
  .s_axi_rvalid(DMA_S_AXI_rvalid),      // output wire s_axi_rvalid
  .s_axi_rready(DMA_S_AXI_rready),      // input wire s_axi_rready


  .m_axi_aclk(firesim_internal_clock),          // input wire m_axi_aclk
  .m_axi_aresetn(rst_firesim_n_sync),    // input wire m_axi_aresetn

  .m_axi_awid(sh_cl_dma_pcis_awid_FIRESIM),          // output wire [5 : 0] m_axi_awid
  .m_axi_awaddr(sh_cl_dma_pcis_awaddr_FIRESIM),      // output wire [63 : 0] m_axi_awaddr
  .m_axi_awlen(sh_cl_dma_pcis_awlen_FIRESIM),        // output wire [7 : 0] m_axi_awlen
  .m_axi_awsize(sh_cl_dma_pcis_awsize_FIRESIM),      // output wire [2 : 0] m_axi_awsize
  .m_axi_awburst(),    // output wire [1 : 0] m_axi_awburst
  .m_axi_awlock(),      // output wire [0 : 0] m_axi_awlock
  .m_axi_awcache(),    // output wire [3 : 0] m_axi_awcache
  .m_axi_awprot(),      // output wire [2 : 0] m_axi_awprot
  .m_axi_awregion(),  // output wire [3 : 0] m_axi_awregion
  .m_axi_awqos(),        // output wire [3 : 0] m_axi_awqos
  .m_axi_awvalid(sh_cl_dma_pcis_awvalid_FIRESIM),    // output wire m_axi_awvalid
  .m_axi_awready(cl_sh_dma_pcis_awready_FIRESIM),    // input wire m_axi_awready

  .m_axi_wdata(sh_cl_dma_pcis_wdata_FIRESIM),        // output wire [511 : 0] m_axi_wdata
  .m_axi_wstrb(sh_cl_dma_pcis_wstrb_FIRESIM),        // output wire [63 : 0] m_axi_wstrb
  .m_axi_wlast(sh_cl_dma_pcis_wlast_FIRESIM),        // output wire m_axi_wlast
  .m_axi_wvalid(sh_cl_dma_pcis_wvalid_FIRESIM),      // output wire m_axi_wvalid
  .m_axi_wready(cl_sh_dma_pcis_wready_FIRESIM),      // input wire m_axi_wready

  .m_axi_bid(cl_sh_dma_pcis_bid_FIRESIM_wide),            // input wire [5 : 0] m_axi_bid
  .m_axi_bresp(cl_sh_dma_pcis_bresp_FIRESIM),        // input wire [1 : 0] m_axi_bresp
  .m_axi_bvalid(cl_sh_dma_pcis_bvalid_FIRESIM),      // input wire m_axi_bvalid
  .m_axi_bready(sh_cl_dma_pcis_bready_FIRESIM),      // output wire m_axi_bready

  .m_axi_arid(sh_cl_dma_pcis_arid_FIRESIM),          // output wire [5 : 0] m_axi_arid
  .m_axi_araddr(sh_cl_dma_pcis_araddr_FIRESIM),      // output wire [63 : 0] m_axi_araddr
  .m_axi_arlen(sh_cl_dma_pcis_arlen_FIRESIM),        // output wire [7 : 0] m_axi_arlen
  .m_axi_arsize(sh_cl_dma_pcis_arsize_FIRESIM),      // output wire [2 : 0] m_axi_arsize
  .m_axi_arburst(),    // output wire [1 : 0] m_axi_arburst
  .m_axi_arlock(),      // output wire [0 : 0] m_axi_arlock
  .m_axi_arcache(),    // output wire [3 : 0] m_axi_arcache
  .m_axi_arprot(),      // output wire [2 : 0] m_axi_arprot
  .m_axi_arregion(),  // output wire [3 : 0] m_axi_arregion
  .m_axi_arqos(),        // output wire [3 : 0] m_axi_arqos
  .m_axi_arvalid(sh_cl_dma_pcis_arvalid_FIRESIM),    // output wire m_axi_arvalid
  .m_axi_arready(cl_sh_dma_pcis_arready_FIRESIM),    // input wire m_axi_arready

  .m_axi_rid(cl_sh_dma_pcis_rid_FIRESIM_wide),            // input wire [5 : 0] m_axi_rid
  .m_axi_rdata(cl_sh_dma_pcis_rdata_FIRESIM),        // input wire [511 : 0] m_axi_rdata
  .m_axi_rresp(cl_sh_dma_pcis_rresp_FIRESIM),        // input wire [1 : 0] m_axi_rresp
  .m_axi_rlast(cl_sh_dma_pcis_rlast_FIRESIM),        // input wire m_axi_rlast
  .m_axi_rvalid(cl_sh_dma_pcis_rvalid_FIRESIM),      // input wire m_axi_rvalid
  .m_axi_rready(sh_cl_dma_pcis_rready_FIRESIM)      // output wire m_axi_rready
);





//----------------------------------------- 
// DDR controller instantiation   
//-----------------------------------------

// Defining local parameters that will instantiate the
// 3 DRAM controllers inside the CL
  
localparam DDR_A_PRESENT = `USE_DDR_CHANNEL_A;

// Define the addition pipeline stag
// needed to close timing for the various
// place where ATG (Automatic Test Generator)
// is defined
   
localparam NUM_CFG_STGS_CL_DDR_ATG = 8;
localparam NUM_CFG_STGS_SH_DDR_ATG = 4;
localparam NUM_CFG_STGS_PCIE_ATG = 4;


// To reduce RTL simulation time, only 8KiB of
// each external DRAM is scrubbed in simulations

`ifdef SIM
   localparam DDR_SCRB_MAX_ADDR = 64'h1FFF;
`else   
   localparam DDR_SCRB_MAX_ADDR = 64'h3FFFFFFFF; //16GB 
`endif
   localparam DDR_SCRB_BURST_LEN_MINUS1 = 15;

`ifdef NO_CL_TST_SCRUBBER
   localparam NO_SCRB_INST = 1;
`else
   localparam NO_SCRB_INST = 0;
`endif   

//-------------------------------------------------------------------------------
//================================================================================
//------------------------------------------------------------------------------

wire [33 : 0] fsimtop_s_0_axi_awaddr_small;
wire [33 : 0] fsimtop_s_0_axi_araddr_small;

wire [15 : 0] fsimtop_s_0_axi_awid;
wire [5 : 0] fsimtop_s_0_axi_awid_short;
assign fsimtop_s_0_axi_awid = {10'b0, fsimtop_s_0_axi_awid_short};

wire [63 : 0] fsimtop_s_0_axi_awaddr;
assign fsimtop_s_0_axi_awaddr = { 30'b0, fsimtop_s_0_axi_awaddr_small[33:0] };
wire [7 : 0] fsimtop_s_0_axi_awlen;
wire [2 : 0] fsimtop_s_0_axi_awsize;
wire [1 : 0] fsimtop_s_0_axi_awburst;
wire [0 : 0] fsimtop_s_0_axi_awlock;
wire [3 : 0] fsimtop_s_0_axi_awcache;
wire [2 : 0] fsimtop_s_0_axi_awprot;
wire [3 : 0] fsimtop_s_0_axi_awregion = 4'b0;
wire [3 : 0] fsimtop_s_0_axi_awqos;
wire fsimtop_s_0_axi_awvalid;
wire fsimtop_s_0_axi_awready;

wire [63 : 0] fsimtop_s_0_axi_wdata;
wire [7 : 0] fsimtop_s_0_axi_wstrb;
wire fsimtop_s_0_axi_wlast;
wire fsimtop_s_0_axi_wvalid;
wire fsimtop_s_0_axi_wready;

wire [15 : 0] fsimtop_s_0_axi_bid;
wire [1 : 0] fsimtop_s_0_axi_bresp;
wire fsimtop_s_0_axi_bvalid;
wire fsimtop_s_0_axi_bready;

wire [15 : 0] fsimtop_s_0_axi_arid;
wire [5 : 0] fsimtop_s_0_axi_arid_short;
assign fsimtop_s_0_axi_arid = {10'b0, fsimtop_s_0_axi_arid_short};

wire [63 : 0] fsimtop_s_0_axi_araddr;
assign fsimtop_s_0_axi_araddr = { 30'b0, fsimtop_s_0_axi_araddr_small[33:0] };
wire [7 : 0] fsimtop_s_0_axi_arlen;
wire [2 : 0] fsimtop_s_0_axi_arsize;
wire [1 : 0] fsimtop_s_0_axi_arburst;
wire [0 : 0] fsimtop_s_0_axi_arlock;
wire [3 : 0] fsimtop_s_0_axi_arcache;
wire [2 : 0] fsimtop_s_0_axi_arprot;
wire [3 : 0] fsimtop_s_0_axi_arregion = 4'b0;
wire [3 : 0] fsimtop_s_0_axi_arqos;
wire fsimtop_s_0_axi_arvalid;
wire fsimtop_s_0_axi_arready;

wire [15 : 0] fsimtop_s_0_axi_rid;
wire [63 : 0] fsimtop_s_0_axi_rdata;
wire [1 : 0] fsimtop_s_0_axi_rresp;
wire fsimtop_s_0_axi_rlast;
wire fsimtop_s_0_axi_rvalid;
wire fsimtop_s_0_axi_rready;


wire [33 : 0] fsimtop_s_1_axi_awaddr_small;
wire [33 : 0] fsimtop_s_1_axi_araddr_small;

wire [15 : 0] fsimtop_s_1_axi_awid;
wire [5 : 0] fsimtop_s_1_axi_awid_short;
assign fsimtop_s_1_axi_awid = {10'b0, fsimtop_s_1_axi_awid_short};

wire [63 : 0] fsimtop_s_1_axi_awaddr;
assign fsimtop_s_1_axi_awaddr = { 30'b0, fsimtop_s_1_axi_awaddr_small[33:0] };
wire [7 : 0] fsimtop_s_1_axi_awlen;
wire [2 : 0] fsimtop_s_1_axi_awsize;
wire [1 : 0] fsimtop_s_1_axi_awburst;
wire [0 : 0] fsimtop_s_1_axi_awlock;
wire [3 : 0] fsimtop_s_1_axi_awcache;
wire [2 : 0] fsimtop_s_1_axi_awprot;
wire [3 : 0] fsimtop_s_1_axi_awregion = 4'b0;
wire [3 : 0] fsimtop_s_1_axi_awqos;
wire fsimtop_s_1_axi_awvalid;
wire fsimtop_s_1_axi_awready;

wire [63 : 0] fsimtop_s_1_axi_wdata;
wire [7 : 0] fsimtop_s_1_axi_wstrb;
wire fsimtop_s_1_axi_wlast;
wire fsimtop_s_1_axi_wvalid;
wire fsimtop_s_1_axi_wready;

wire [15 : 0] fsimtop_s_1_axi_bid;
wire [1 : 0] fsimtop_s_1_axi_bresp;
wire fsimtop_s_1_axi_bvalid;
wire fsimtop_s_1_axi_bready;

wire [15 : 0] fsimtop_s_1_axi_arid;
wire [5 : 0] fsimtop_s_1_axi_arid_short;
assign fsimtop_s_1_axi_arid = {10'b0, fsimtop_s_1_axi_arid_short};

wire [63 : 0] fsimtop_s_1_axi_araddr;
assign fsimtop_s_1_axi_araddr = { 30'b0, fsimtop_s_1_axi_araddr_small[33:0] };
wire [7 : 0] fsimtop_s_1_axi_arlen;
wire [2 : 0] fsimtop_s_1_axi_arsize;
wire [1 : 0] fsimtop_s_1_axi_arburst;
wire [0 : 0] fsimtop_s_1_axi_arlock;
wire [3 : 0] fsimtop_s_1_axi_arcache;
wire [2 : 0] fsimtop_s_1_axi_arprot;
wire [3 : 0] fsimtop_s_1_axi_arregion = 4'b0;
wire [3 : 0] fsimtop_s_1_axi_arqos;
wire fsimtop_s_1_axi_arvalid;
wire fsimtop_s_1_axi_arready;

wire [15 : 0] fsimtop_s_1_axi_rid;
wire [63 : 0] fsimtop_s_1_axi_rdata;
wire [1 : 0] fsimtop_s_1_axi_rresp;
wire fsimtop_s_1_axi_rlast;
wire fsimtop_s_1_axi_rvalid;
wire fsimtop_s_1_axi_rready;



  F1Shim firesim_top (
   .clock(firesim_internal_clock),
   .reset(!rst_firesim_n_sync),
   .io_master_aw_ready(ocl_sh_awready_q),
   .io_master_aw_valid(sh_ocl_awvalid_q),
   .io_master_aw_bits_addr(sh_ocl_awaddr_q[24:0]),
   .io_master_aw_bits_len(8'h0),
   .io_master_aw_bits_size(3'h2),
   .io_master_aw_bits_burst(2'h1),
   .io_master_aw_bits_lock(1'h0),
   .io_master_aw_bits_cache(4'h0),
   .io_master_aw_bits_prot(3'h0), //unused? (could connect?)
   .io_master_aw_bits_qos(4'h0),
   .io_master_aw_bits_region(4'h0),
   .io_master_aw_bits_id(12'h0),
   .io_master_aw_bits_user(1'h0),
   .io_master_w_ready(ocl_sh_wready_q),
   .io_master_w_valid(sh_ocl_wvalid_q),
   .io_master_w_bits_data(sh_ocl_wdata_q),
   .io_master_w_bits_last(1'h1),
   .io_master_w_bits_id(12'h0),
   .io_master_w_bits_strb(sh_ocl_wstrb_q), //OR 8'hff
   .io_master_w_bits_user(1'h0),
   .io_master_b_ready(sh_ocl_bready_q),
   .io_master_b_valid(ocl_sh_bvalid_q),
   .io_master_b_bits_resp(ocl_sh_bresp_q),
   .io_master_b_bits_id(),      // UNUSED at top level
   .io_master_b_bits_user(),    // UNUSED at top level
   .io_master_ar_ready(ocl_sh_arready_q),
   .io_master_ar_valid(sh_ocl_arvalid_q),
   .io_master_ar_bits_addr(sh_ocl_araddr_q[24:0]),
   .io_master_ar_bits_len(8'h0),
   .io_master_ar_bits_size(3'h2),
   .io_master_ar_bits_burst(2'h1),
   .io_master_ar_bits_lock(1'h0),
   .io_master_ar_bits_cache(4'h0),
   .io_master_ar_bits_prot(3'h0),
   .io_master_ar_bits_qos(4'h0),
   .io_master_ar_bits_region(4'h0),
   .io_master_ar_bits_id(12'h0),
   .io_master_ar_bits_user(1'h0),
   .io_master_r_ready(sh_ocl_rready_q),
   .io_master_r_valid(ocl_sh_rvalid_q),
   .io_master_r_bits_resp(ocl_sh_rresp_q),
   .io_master_r_bits_data(ocl_sh_rdata_q),
   .io_master_r_bits_last(), //UNUSED at top level
   .io_master_r_bits_id(),      // UNUSED at top level
   .io_master_r_bits_user(),    // UNUSED at top level

    // special NIC master interface
   .io_pcis_aw_ready(cl_sh_dma_pcis_awready_FIRESIM),
   .io_pcis_aw_valid(sh_cl_dma_pcis_awvalid_FIRESIM),
   .io_pcis_aw_bits_addr(sh_cl_dma_pcis_awaddr_FIRESIM),
   .io_pcis_aw_bits_len(sh_cl_dma_pcis_awlen_FIRESIM),
   .io_pcis_aw_bits_size(sh_cl_dma_pcis_awsize_FIRESIM),
   .io_pcis_aw_bits_burst(2'h1),
   .io_pcis_aw_bits_lock(1'h0),
   .io_pcis_aw_bits_cache(4'h0),
   .io_pcis_aw_bits_prot(3'h0), //unused? (could connect?)
   .io_pcis_aw_bits_qos(4'h0),
   .io_pcis_aw_bits_region(4'h0),
   .io_pcis_aw_bits_id(sh_cl_dma_pcis_awid_FIRESIM),
   .io_pcis_aw_bits_user(1'h0),
   .io_pcis_w_ready(cl_sh_dma_pcis_wready_FIRESIM),
   .io_pcis_w_valid(sh_cl_dma_pcis_wvalid_FIRESIM),
   .io_pcis_w_bits_data(sh_cl_dma_pcis_wdata_FIRESIM),
   .io_pcis_w_bits_last(sh_cl_dma_pcis_wlast_FIRESIM),
   .io_pcis_w_bits_id(6'h0),
   .io_pcis_w_bits_strb(sh_cl_dma_pcis_wstrb_FIRESIM),
   .io_pcis_w_bits_user(1'h0),
   .io_pcis_b_ready(sh_cl_dma_pcis_bready_FIRESIM),
   .io_pcis_b_valid(cl_sh_dma_pcis_bvalid_FIRESIM),
   .io_pcis_b_bits_resp(cl_sh_dma_pcis_bresp_FIRESIM),
   .io_pcis_b_bits_id(cl_sh_dma_pcis_bid_FIRESIM),
   .io_pcis_b_bits_user(),    // UNUSED at top level
   .io_pcis_ar_ready(cl_sh_dma_pcis_arready_FIRESIM),
   .io_pcis_ar_valid(sh_cl_dma_pcis_arvalid_FIRESIM),
   .io_pcis_ar_bits_addr(sh_cl_dma_pcis_araddr_FIRESIM),
   .io_pcis_ar_bits_len(sh_cl_dma_pcis_arlen_FIRESIM),
   .io_pcis_ar_bits_size(sh_cl_dma_pcis_arsize_FIRESIM),
   .io_pcis_ar_bits_burst(2'h1),
   .io_pcis_ar_bits_lock(1'h0),
   .io_pcis_ar_bits_cache(4'h0),
   .io_pcis_ar_bits_prot(3'h0),
   .io_pcis_ar_bits_qos(4'h0),
   .io_pcis_ar_bits_region(4'h0),
   .io_pcis_ar_bits_id(sh_cl_dma_pcis_arid_FIRESIM),
   .io_pcis_ar_bits_user(1'h0),
   .io_pcis_r_ready(sh_cl_dma_pcis_rready_FIRESIM),
   .io_pcis_r_valid(cl_sh_dma_pcis_rvalid_FIRESIM),
   .io_pcis_r_bits_resp(cl_sh_dma_pcis_rresp_FIRESIM),
   .io_pcis_r_bits_data(cl_sh_dma_pcis_rdata_FIRESIM),
   .io_pcis_r_bits_last(cl_sh_dma_pcis_rlast_FIRESIM),
   .io_pcis_r_bits_id(cl_sh_dma_pcis_rid_FIRESIM),
   .io_pcis_r_bits_user(),    // UNUSED at top level

   .io_slave_0_aw_ready(fsimtop_s_0_axi_awready),
   .io_slave_0_aw_valid(fsimtop_s_0_axi_awvalid),
   .io_slave_0_aw_bits_addr(fsimtop_s_0_axi_awaddr_small),
   .io_slave_0_aw_bits_len(fsimtop_s_0_axi_awlen),
   .io_slave_0_aw_bits_size(fsimtop_s_0_axi_awsize),
   .io_slave_0_aw_bits_burst(fsimtop_s_0_axi_awburst), // not available on DDR IF
   .io_slave_0_aw_bits_lock(fsimtop_s_0_axi_awlock), // not available on DDR IF
   .io_slave_0_aw_bits_cache(fsimtop_s_0_axi_awcache), // not available on DDR IF
   .io_slave_0_aw_bits_prot(fsimtop_s_0_axi_awprot), // not available on DDR IF
   .io_slave_0_aw_bits_qos(fsimtop_s_0_axi_awqos), // not available on DDR IF
   .io_slave_0_aw_bits_id(fsimtop_s_0_axi_awid_short),

   .io_slave_0_w_ready(fsimtop_s_0_axi_wready),
   .io_slave_0_w_valid(fsimtop_s_0_axi_wvalid),
   .io_slave_0_w_bits_data(fsimtop_s_0_axi_wdata),
   .io_slave_0_w_bits_last(fsimtop_s_0_axi_wlast),
   .io_slave_0_w_bits_strb(fsimtop_s_0_axi_wstrb),

   .io_slave_0_b_ready(fsimtop_s_0_axi_bready),
   .io_slave_0_b_valid(fsimtop_s_0_axi_bvalid),
   .io_slave_0_b_bits_resp(fsimtop_s_0_axi_bresp),
   .io_slave_0_b_bits_id(fsimtop_s_0_axi_bid),

   .io_slave_0_ar_ready(fsimtop_s_0_axi_arready),
   .io_slave_0_ar_valid(fsimtop_s_0_axi_arvalid),
   .io_slave_0_ar_bits_addr(fsimtop_s_0_axi_araddr_small),
   .io_slave_0_ar_bits_len(fsimtop_s_0_axi_arlen),
   .io_slave_0_ar_bits_size(fsimtop_s_0_axi_arsize),
   .io_slave_0_ar_bits_burst(fsimtop_s_0_axi_arburst), // not available on DDR IF
   .io_slave_0_ar_bits_lock(fsimtop_s_0_axi_arlock), // not available on DDR IF
   .io_slave_0_ar_bits_cache(fsimtop_s_0_axi_arcache), // not available on DDR IF
   .io_slave_0_ar_bits_prot(fsimtop_s_0_axi_arprot), // not available on DDR IF
   .io_slave_0_ar_bits_qos(fsimtop_s_0_axi_arqos), // not available on DDR IF
   .io_slave_0_ar_bits_id(fsimtop_s_0_axi_arid_short), // not available on DDR IF

   .io_slave_0_r_ready(fsimtop_s_0_axi_rready),
   .io_slave_0_r_valid(fsimtop_s_0_axi_rvalid),
   .io_slave_0_r_bits_resp(fsimtop_s_0_axi_rresp),
   .io_slave_0_r_bits_data(fsimtop_s_0_axi_rdata),
   .io_slave_0_r_bits_last(fsimtop_s_0_axi_rlast),
   .io_slave_0_r_bits_id(fsimtop_s_0_axi_rid),

   .io_slave_1_aw_ready(fsimtop_s_1_axi_awready),
   .io_slave_1_aw_valid(fsimtop_s_1_axi_awvalid),
   .io_slave_1_aw_bits_addr(fsimtop_s_1_axi_awaddr_small),
   .io_slave_1_aw_bits_len(fsimtop_s_1_axi_awlen),
   .io_slave_1_aw_bits_size(fsimtop_s_1_axi_awsize),
   .io_slave_1_aw_bits_burst(fsimtop_s_1_axi_awburst), // not available on DDR IF
   .io_slave_1_aw_bits_lock(fsimtop_s_1_axi_awlock), // not available on DDR IF
   .io_slave_1_aw_bits_cache(fsimtop_s_1_axi_awcache), // not available on DDR IF
   .io_slave_1_aw_bits_prot(fsimtop_s_1_axi_awprot), // not available on DDR IF
   .io_slave_1_aw_bits_qos(fsimtop_s_1_axi_awqos), // not available on DDR IF
   .io_slave_1_aw_bits_id(fsimtop_s_1_axi_awid_short),

   .io_slave_1_w_ready(fsimtop_s_1_axi_wready),
   .io_slave_1_w_valid(fsimtop_s_1_axi_wvalid),
   .io_slave_1_w_bits_data(fsimtop_s_1_axi_wdata),
   .io_slave_1_w_bits_last(fsimtop_s_1_axi_wlast),
   .io_slave_1_w_bits_strb(fsimtop_s_1_axi_wstrb),

   .io_slave_1_b_ready(fsimtop_s_1_axi_bready),
   .io_slave_1_b_valid(fsimtop_s_1_axi_bvalid),
   .io_slave_1_b_bits_resp(fsimtop_s_1_axi_bresp),
   .io_slave_1_b_bits_id(fsimtop_s_1_axi_bid),

   .io_slave_1_ar_ready(fsimtop_s_1_axi_arready),
   .io_slave_1_ar_valid(fsimtop_s_1_axi_arvalid),
   .io_slave_1_ar_bits_addr(fsimtop_s_1_axi_araddr_small),
   .io_slave_1_ar_bits_len(fsimtop_s_1_axi_arlen),
   .io_slave_1_ar_bits_size(fsimtop_s_1_axi_arsize),
   .io_slave_1_ar_bits_burst(fsimtop_s_1_axi_arburst), // not available on DDR IF
   .io_slave_1_ar_bits_lock(fsimtop_s_1_axi_arlock), // not available on DDR IF
   .io_slave_1_ar_bits_cache(fsimtop_s_1_axi_arcache), // not available on DDR IF
   .io_slave_1_ar_bits_prot(fsimtop_s_1_axi_arprot), // not available on DDR IF
   .io_slave_1_ar_bits_qos(fsimtop_s_1_axi_arqos), // not available on DDR IF
   .io_slave_1_ar_bits_id(fsimtop_s_1_axi_arid_short), // not available on DDR IF

   .io_slave_1_r_ready(fsimtop_s_1_axi_rready),
   .io_slave_1_r_valid(fsimtop_s_1_axi_rvalid),
   .io_slave_1_r_bits_resp(fsimtop_s_1_axi_rresp),
   .io_slave_1_r_bits_data(fsimtop_s_1_axi_rdata),
   .io_slave_1_r_bits_last(fsimtop_s_1_axi_rlast),
   .io_slave_1_r_bits_id(fsimtop_s_1_axi_rid)
);

//****************DDR CHANNEL C****************************

wire [15 : 0] clock_converted_axi_0_awid;
wire [63 : 0] clock_converted_axi_0_awaddr;
wire [7 : 0]  clock_converted_axi_0_awlen;
wire [2 : 0]  clock_converted_axi_0_awsize;
wire [1 : 0]  clock_converted_axi_0_awburst;
wire [0 : 0]  clock_converted_axi_0_awlock;
wire [3 : 0]  clock_converted_axi_0_awcache;
wire [2 : 0]  clock_converted_axi_0_awprot;
wire [3 : 0]  clock_converted_axi_0_awregion;
wire [3 : 0]  clock_converted_axi_0_awqos;
wire          clock_converted_axi_0_awvalid;
wire          clock_converted_axi_0_awready;

wire [63 : 0] clock_converted_axi_0_wdata;
wire [7 : 0]  clock_converted_axi_0_wstrb;
wire          clock_converted_axi_0_wlast;
wire          clock_converted_axi_0_wvalid;
wire          clock_converted_axi_0_wready;

wire [15 : 0] clock_converted_axi_0_bid;
wire [1 : 0]  clock_converted_axi_0_bresp;
wire          clock_converted_axi_0_bvalid;
wire          clock_converted_axi_0_bready;

wire [15 : 0] clock_converted_axi_0_arid;
wire [63 : 0] clock_converted_axi_0_araddr;
wire [7 : 0]  clock_converted_axi_0_arlen;
wire [2 : 0]  clock_converted_axi_0_arsize;
wire [1 : 0]  clock_converted_axi_0_arburst;
wire [0 : 0]  clock_converted_axi_0_arlock;
wire [3 : 0]  clock_converted_axi_0_arcache;
wire [2 : 0]  clock_converted_axi_0_arprot;
wire [3 : 0]  clock_converted_axi_0_arregion;
wire [3 : 0]  clock_converted_axi_0_arqos;
wire          clock_converted_axi_0_arvalid;
wire          clock_converted_axi_0_arready;

wire [15 : 0] clock_converted_axi_0_rid;
wire [63 : 0] clock_converted_axi_0_rdata;
wire [1 : 0]  clock_converted_axi_0_rresp;
wire          clock_converted_axi_0_rlast;
wire          clock_converted_axi_0_rvalid;
wire          clock_converted_axi_0_rready;

axi_clock_converter_dramslim clock_convert_dramslim_0 (
  .s_axi_aclk(firesim_internal_clock),          // input wire s_axi_aclk
  .s_axi_aresetn(rst_firesim_n_sync),    // input wire s_axi_aresetn

  .s_axi_awid(fsimtop_s_0_axi_awid),          // input wire [15 : 0] s_axi_awid
  .s_axi_awaddr(fsimtop_s_0_axi_awaddr),      // input wire [63 : 0] s_axi_awaddr
  .s_axi_awlen(fsimtop_s_0_axi_awlen),        // input wire [7 : 0] s_axi_awlen
  .s_axi_awsize(fsimtop_s_0_axi_awsize),      // input wire [2 : 0] s_axi_awsize
  .s_axi_awburst(fsimtop_s_0_axi_awburst),    // input wire [1 : 0] s_axi_awburst
  .s_axi_awlock(fsimtop_s_0_axi_awlock),      // input wire [0 : 0] s_axi_awlock
  // CACHE = xx1x indicates the transcation is modifiable and
  // that the converter should pack narrow writes into wider ones
  .s_axi_awcache(4'h2),    // input wire [3 : 0] s_axi_awcache
  .s_axi_awprot(fsimtop_s_0_axi_awprot),      // input wire [2 : 0] s_axi_awprot
  .s_axi_awregion(fsimtop_s_0_axi_awregion),  // input wire [3 : 0] s_axi_awregion
  .s_axi_awqos(fsimtop_s_0_axi_awqos),        // input wire [3 : 0] s_axi_awqos
  .s_axi_awvalid(fsimtop_s_0_axi_awvalid),    // input wire s_axi_awvalid
  .s_axi_awready(fsimtop_s_0_axi_awready),    // output wire s_axi_awready

  .s_axi_wdata(fsimtop_s_0_axi_wdata),        // input wire [63 : 0] s_axi_wdata
  .s_axi_wstrb(fsimtop_s_0_axi_wstrb),        // input wire [7 : 0] s_axi_wstrb
  .s_axi_wlast(fsimtop_s_0_axi_wlast),        // input wire s_axi_wlast
  .s_axi_wvalid(fsimtop_s_0_axi_wvalid),      // input wire s_axi_wvalid
  .s_axi_wready(fsimtop_s_0_axi_wready),      // output wire s_axi_wready

  .s_axi_bid(fsimtop_s_0_axi_bid),            // output wire [15 : 0] s_axi_bid
  .s_axi_bresp(fsimtop_s_0_axi_bresp),        // output wire [1 : 0] s_axi_bresp
  .s_axi_bvalid(fsimtop_s_0_axi_bvalid),      // output wire s_axi_bvalid
  .s_axi_bready(fsimtop_s_0_axi_bready),      // input wire s_axi_bready

  .s_axi_arid(fsimtop_s_0_axi_arid),          // input wire [15 : 0] s_axi_arid
  .s_axi_araddr(fsimtop_s_0_axi_araddr),      // input wire [63 : 0] s_axi_araddr
  .s_axi_arlen(fsimtop_s_0_axi_arlen),        // input wire [7 : 0] s_axi_arlen
  .s_axi_arsize(fsimtop_s_0_axi_arsize),      // input wire [2 : 0] s_axi_arsize
  .s_axi_arburst(fsimtop_s_0_axi_arburst),    // input wire [1 : 0] s_axi_arburst
  .s_axi_arlock(fsimtop_s_0_axi_arlock),      // input wire [0 : 0] s_axi_arlock
  // CACHE = xx1x indicates the transcation is modifiable and
  // that the converter should pack narrow reads into wider ones
  .s_axi_arcache(4'h2),                     // input wire [3 : 0] s_axi_arcache
  .s_axi_arprot(fsimtop_s_0_axi_arprot),      // input wire [2 : 0] s_axi_arprot
  .s_axi_arregion(fsimtop_s_0_axi_arregion),  // input wire [3 : 0] s_axi_arregion
  .s_axi_arqos(fsimtop_s_0_axi_arqos),        // input wire [3 : 0] s_axi_arqos
  .s_axi_arvalid(fsimtop_s_0_axi_arvalid),    // input wire s_axi_arvalid
  .s_axi_arready(fsimtop_s_0_axi_arready),    // output wire s_axi_arready

  .s_axi_rid(fsimtop_s_0_axi_rid),            // output wire [15 : 0] s_axi_rid
  .s_axi_rdata(fsimtop_s_0_axi_rdata),        // output wire [63 : 0] s_axi_rdata
  .s_axi_rresp(fsimtop_s_0_axi_rresp),        // output wire [1 : 0] s_axi_rresp
  .s_axi_rlast(fsimtop_s_0_axi_rlast),        // output wire s_axi_rlast
  .s_axi_rvalid(fsimtop_s_0_axi_rvalid),      // output wire s_axi_rvalid
  .s_axi_rready(fsimtop_s_0_axi_rready),      // input wire s_axi_rready

  .m_axi_aclk(clk),          // input wire m_axi_aclk
  .m_axi_aresetn(rst_main_n_sync),    // input wire m_axi_aresetn

  .m_axi_awid(clock_converted_axi_0_awid),          // output wire [15 : 0] m_axi_awid
  .m_axi_awaddr(clock_converted_axi_0_awaddr),      // output wire [63 : 0] m_axi_awaddr
  .m_axi_awlen(clock_converted_axi_0_awlen),        // output wire [7 : 0] m_axi_awlen
  .m_axi_awsize(clock_converted_axi_0_awsize),      // output wire [2 : 0] m_axi_awsize
  .m_axi_awburst(clock_converted_axi_0_awburst),    // output wire [1 : 0] m_axi_awburst
  .m_axi_awlock(clock_converted_axi_0_awlock),      // output wire [0 : 0] m_axi_awlock
  .m_axi_awcache(clock_converted_axi_0_awcache),    // output wire [3 : 0] m_axi_awcache
  .m_axi_awprot(clock_converted_axi_0_awprot),      // output wire [2 : 0] m_axi_awprot
  .m_axi_awregion(clock_converted_axi_0_awregion),  // output wire [3 : 0] m_axi_awregion
  .m_axi_awqos(clock_converted_axi_0_awqos),        // output wire [3 : 0] m_axi_awqos
  .m_axi_awvalid(clock_converted_axi_0_awvalid),    // output wire m_axi_awvalid
  .m_axi_awready(clock_converted_axi_0_awready),    // input wire m_axi_awready

  .m_axi_wdata(clock_converted_axi_0_wdata),        // output wire [511 : 0] m_axi_wdata
  .m_axi_wstrb(clock_converted_axi_0_wstrb),        // output wire [63 : 0] m_axi_wstrb
  .m_axi_wlast(clock_converted_axi_0_wlast),        // output wire m_axi_wlast
  .m_axi_wvalid(clock_converted_axi_0_wvalid),      // output wire m_axi_wvalid
  .m_axi_wready(clock_converted_axi_0_wready),      // input wire m_axi_wready

  .m_axi_bid(clock_converted_axi_0_bid),            // input wire [15 : 0] m_axi_bid
  .m_axi_bresp(clock_converted_axi_0_bresp),        // input wire [1 : 0] m_axi_bresp
  .m_axi_bvalid(clock_converted_axi_0_bvalid),      // input wire m_axi_bvalid
  .m_axi_bready(clock_converted_axi_0_bready),      // output wire m_axi_bready

  .m_axi_arid(clock_converted_axi_0_arid),          // output wire [15 : 0] m_axi_arid
  .m_axi_araddr(clock_converted_axi_0_araddr),      // output wire [63 : 0] m_axi_araddr
  .m_axi_arlen(clock_converted_axi_0_arlen),        // output wire [7 : 0] m_axi_arlen
  .m_axi_arsize(clock_converted_axi_0_arsize),      // output wire [2 : 0] m_axi_arsize
  .m_axi_arburst(clock_converted_axi_0_arburst),    // output wire [1 : 0] m_axi_arburst
  .m_axi_arlock(clock_converted_axi_0_arlock),      // output wire [0 : 0] m_axi_arlock
  .m_axi_arcache(clock_converted_axi_0_arcache),    // output wire [3 : 0] m_axi_arcache
  .m_axi_arprot(clock_converted_axi_0_arprot),      // output wire [2 : 0] m_axi_arprot
  .m_axi_arregion(clock_converted_axi_0_arregion),  // output wire [3 : 0] m_axi_arregion
  .m_axi_arqos(clock_converted_axi_0_arqos),        // output wire [3 : 0] m_axi_arqos
  .m_axi_arvalid(clock_converted_axi_0_arvalid),    // output wire m_axi_arvalid
  .m_axi_arready(clock_converted_axi_0_arready),    // input wire m_axi_arready

  .m_axi_rid(clock_converted_axi_0_rid),            // input wire [15 : 0] m_axi_rid
  .m_axi_rdata(clock_converted_axi_0_rdata),        // input wire [511 : 0] m_axi_rdata
  .m_axi_rresp(clock_converted_axi_0_rresp),        // input wire [1 : 0] m_axi_rresp
  .m_axi_rlast(clock_converted_axi_0_rlast),        // input wire m_axi_rlast
  .m_axi_rvalid(clock_converted_axi_0_rvalid),      // input wire m_axi_rvalid
  .m_axi_rready(clock_converted_axi_0_rready)      // output wire m_axi_rready
);

/* steps to move:
 * 1) copy clock converter's M interfaces to dwidth converter's M interfaces: DONE
 * 2) create clock_converted_* signals for clock M to width adapt S: DONE
 * 3) add asserts on arsize and awsize to confirm that they're always b110
*/

assign DDRA_M_AXI_awid = 16'b0; // dwidth convert has no awid for some reason...
assign DDRA_M_AXI_arid = 16'b0; // dwidth convert has no arid for some reason...
// unused: sh_cl_ddr_bid
// unused: sh_cl_ddr_rid

axi_dwidth_converter_0 dwidth_adapt_64bits_512bits_0 (
  .s_axi_aclk(clk),          // input wire s_axi_aclk
  .s_axi_aresetn(rst_main_n_sync),    // input wire s_axi_aresetn

  .s_axi_awid(clock_converted_axi_0_awid),          // input wire [15 : 0] s_axi_awid
  .s_axi_awaddr(clock_converted_axi_0_awaddr),      // input wire [63 : 0] s_axi_awaddr
  .s_axi_awlen(clock_converted_axi_0_awlen),        // input wire [7 : 0] s_axi_awlen
  .s_axi_awsize(clock_converted_axi_0_awsize),      // input wire [2 : 0] s_axi_awsize
  .s_axi_awburst(clock_converted_axi_0_awburst),    // input wire [1 : 0] s_axi_awburst
  .s_axi_awlock(clock_converted_axi_0_awlock),      // input wire [0 : 0] s_axi_awlock
  .s_axi_awcache(clock_converted_axi_0_awcache),    // input wire [3 : 0] s_axi_awcache
  .s_axi_awprot(clock_converted_axi_0_awprot),      // input wire [2 : 0] s_axi_awprot
  .s_axi_awregion(clock_converted_axi_0_awregion),  // input wire [3 : 0] s_axi_awregion
  .s_axi_awqos(clock_converted_axi_0_awqos),        // input wire [3 : 0] s_axi_awqos
  .s_axi_awvalid(clock_converted_axi_0_awvalid),    // input wire s_axi_awvalid
  .s_axi_awready(clock_converted_axi_0_awready),    // output wire s_axi_awready

  .s_axi_wdata(clock_converted_axi_0_wdata),        // input wire [63 : 0] s_axi_wdata
  .s_axi_wstrb(clock_converted_axi_0_wstrb),        // input wire [7 : 0] s_axi_wstrb
  .s_axi_wlast(clock_converted_axi_0_wlast),        // input wire s_axi_wlast
  .s_axi_wvalid(clock_converted_axi_0_wvalid),      // input wire s_axi_wvalid
  .s_axi_wready(clock_converted_axi_0_wready),      // output wire s_axi_wready

  .s_axi_bid(clock_converted_axi_0_bid),            // output wire [15 : 0] s_axi_bid
  .s_axi_bresp(clock_converted_axi_0_bresp),        // output wire [1 : 0] s_axi_bresp
  .s_axi_bvalid(clock_converted_axi_0_bvalid),      // output wire s_axi_bvalid
  .s_axi_bready(clock_converted_axi_0_bready),      // input wire s_axi_bready

  .s_axi_arid(clock_converted_axi_0_arid),          // input wire [15 : 0] s_axi_arid
  .s_axi_araddr(clock_converted_axi_0_araddr),      // input wire [63 : 0] s_axi_araddr
  .s_axi_arlen(clock_converted_axi_0_arlen),        // input wire [7 : 0] s_axi_arlen
  .s_axi_arsize(clock_converted_axi_0_arsize),      // input wire [2 : 0] s_axi_arsize
  .s_axi_arburst(clock_converted_axi_0_arburst),    // input wire [1 : 0] s_axi_arburst
  .s_axi_arlock(clock_converted_axi_0_arlock),      // input wire [0 : 0] s_axi_arlock
  .s_axi_arcache(clock_converted_axi_0_arcache),    // input wire [3 : 0] s_axi_arcache
  .s_axi_arprot(clock_converted_axi_0_arprot),      // input wire [2 : 0] s_axi_arprot
  .s_axi_arregion(clock_converted_axi_0_arregion),  // input wire [3 : 0] s_axi_arregion
  .s_axi_arqos(clock_converted_axi_0_arqos),        // input wire [3 : 0] s_axi_arqos
  .s_axi_arvalid(clock_converted_axi_0_arvalid),    // input wire s_axi_arvalid
  .s_axi_arready(clock_converted_axi_0_arready),    // output wire s_axi_arready

  .s_axi_rid(clock_converted_axi_0_rid),            // output wire [15 : 0] s_axi_rid
  .s_axi_rdata(clock_converted_axi_0_rdata),        // output wire [63 : 0] s_axi_rdata
  .s_axi_rresp(clock_converted_axi_0_rresp),        // output wire [1 : 0] s_axi_rresp
  .s_axi_rlast(clock_converted_axi_0_rlast),        // output wire s_axi_rlast
  .s_axi_rvalid(clock_converted_axi_0_rvalid),      // output wire s_axi_rvalid
  .s_axi_rready(clock_converted_axi_0_rready),      // input wire s_axi_rready


  .m_axi_awaddr(DDRA_M_AXI_awaddr),      // output wire [63 : 0] m_axi_awaddr
  .m_axi_awlen(DDRA_M_AXI_awlen),        // output wire [7 : 0] m_axi_awlen
  .m_axi_awsize(DDRA_M_AXI_awsize),      // output wire [2 : 0] m_axi_awsize
  .m_axi_awburst(DDRA_M_AXI_awburst),    // output wire [1 : 0] m_axi_awburst
  .m_axi_awlock(DDRA_M_AXI_awlock),      // output wire [0 : 0] m_axi_awlock
  .m_axi_awcache(DDRA_M_AXI_awcache),    // output wire [3 : 0] m_axi_awcache
  .m_axi_awprot(DDRA_M_AXI_awprot),      // output wire [2 : 0] m_axi_awprot
  .m_axi_awregion(DDRA_M_AXI_awregion),  // output wire [3 : 0] m_axi_awregion
  .m_axi_awqos(DDRA_M_AXI_awqos),        // output wire [3 : 0] m_axi_awqos
  .m_axi_awvalid(DDRA_M_AXI_awvalid),    // output wire m_axi_awvalid
  .m_axi_awready(DDRA_M_AXI_awready),    // input wire m_axi_awready

  .m_axi_wdata(DDRA_M_AXI_wdata),        // output wire [511 : 0] m_axi_wdata
  .m_axi_wstrb(DDRA_M_AXI_wstrb),        // output wire [63 : 0] m_axi_wstrb
  .m_axi_wlast(DDRA_M_AXI_wlast),        // output wire m_axi_wlast
  .m_axi_wvalid(DDRA_M_AXI_wvalid),      // output wire m_axi_wvalid
  .m_axi_wready(DDRA_M_AXI_wready),      // input wire m_axi_wready

  .m_axi_bresp(DDRA_M_AXI_bresp),        // input wire [1 : 0] m_axi_bresp
  .m_axi_bvalid(DDRA_M_AXI_bvalid),      // input wire m_axi_bvalid
  .m_axi_bready(DDRA_M_AXI_bready),      // output wire m_axi_bready

  .m_axi_araddr(DDRA_M_AXI_araddr),      // output wire [63 : 0] m_axi_araddr
  .m_axi_arlen(DDRA_M_AXI_arlen),        // output wire [7 : 0] m_axi_arlen
  .m_axi_arsize(DDRA_M_AXI_arsize),      // output wire [2 : 0] m_axi_arsize
  .m_axi_arburst(DDRA_M_AXI_arburst),    // output wire [1 : 0] m_axi_arburst
  .m_axi_arlock(DDRA_M_AXI_arlock),      // output wire [0 : 0] m_axi_arlock
  .m_axi_arcache(DDRA_M_AXI_arcache),    // output wire [3 : 0] m_axi_arcache
  .m_axi_arprot(DDRA_M_AXI_arprot),      // output wire [2 : 0] m_axi_arprot
  .m_axi_arregion(DDRA_M_AXI_arregion),  // output wire [3 : 0] m_axi_arregion
  .m_axi_arqos(DDRA_M_AXI_arqos),        // output wire [3 : 0] m_axi_arqos
  .m_axi_arvalid(DDRA_M_AXI_arvalid),    // output wire m_axi_arvalid
  .m_axi_arready(DDRA_M_AXI_arready),    // input wire m_axi_arready

  .m_axi_rdata(DDRA_M_AXI_rdata),        // input wire [511 : 0] m_axi_rdata
  .m_axi_rresp(DDRA_M_AXI_rresp),        // input wire [1 : 0] m_axi_rresp
  .m_axi_rlast(DDRA_M_AXI_rlast),        // input wire m_axi_rlast
  .m_axi_rvalid(DDRA_M_AXI_rvalid),      // input wire m_axi_rvalid
  .m_axi_rready(DDRA_M_AXI_rready)      // output wire m_axi_rready
);



//****************DDR CHANNEL A****************************
generate
    if (DDR_A_PRESENT) begin
        wire [15 : 0] clock_converted_axi_1_awid;
        wire [63 : 0] clock_converted_axi_1_awaddr;
        wire [7 : 0]  clock_converted_axi_1_awlen;
        wire [2 : 0]  clock_converted_axi_1_awsize;
        wire [1 : 0]  clock_converted_axi_1_awburst;
        wire [0 : 0]  clock_converted_axi_1_awlock;
        wire [3 : 0]  clock_converted_axi_1_awcache;
        wire [2 : 0]  clock_converted_axi_1_awprot;
        wire [3 : 0]  clock_converted_axi_1_awregion;
        wire [3 : 0]  clock_converted_axi_1_awqos;
        wire          clock_converted_axi_1_awvalid;
        wire          clock_converted_axi_1_awready;

        wire [63 : 0] clock_converted_axi_1_wdata;
        wire [7 : 0]  clock_converted_axi_1_wstrb;
        wire          clock_converted_axi_1_wlast;
        wire          clock_converted_axi_1_wvalid;
        wire          clock_converted_axi_1_wready;

        wire [15 : 0] clock_converted_axi_1_bid;
        wire [1 : 0]  clock_converted_axi_1_bresp;
        wire          clock_converted_axi_1_bvalid;
        wire          clock_converted_axi_1_bready;

        wire [15 : 0] clock_converted_axi_1_arid;
        wire [63 : 0] clock_converted_axi_1_araddr;
        wire [7 : 0]  clock_converted_axi_1_arlen;
        wire [2 : 0]  clock_converted_axi_1_arsize;
        wire [1 : 0]  clock_converted_axi_1_arburst;
        wire [0 : 0]  clock_converted_axi_1_arlock;
        wire [3 : 0]  clock_converted_axi_1_arcache;
        wire [2 : 0]  clock_converted_axi_1_arprot;
        wire [3 : 0]  clock_converted_axi_1_arregion;
        wire [3 : 0]  clock_converted_axi_1_arqos;
        wire          clock_converted_axi_1_arvalid;
        wire          clock_converted_axi_1_arready;

        wire [15 : 0] clock_converted_axi_1_rid;
        wire [63 : 0] clock_converted_axi_1_rdata;
        wire [1 : 0]  clock_converted_axi_1_rresp;
        wire          clock_converted_axi_1_rlast;
        wire          clock_converted_axi_1_rvalid;
        wire          clock_converted_axi_1_rready;

        axi_clock_converter_dramslim clock_convert_dramslim_1 (
          .s_axi_aclk(firesim_internal_clock),          // input wire s_axi_aclk
          .s_axi_aresetn(rst_firesim_n_sync),    // input wire s_axi_aresetn

          .s_axi_awid(fsimtop_s_1_axi_awid),          // input wire [15 : 0] s_axi_awid
          .s_axi_awaddr(fsimtop_s_1_axi_awaddr),      // input wire [63 : 0] s_axi_awaddr
          .s_axi_awlen(fsimtop_s_1_axi_awlen),        // input wire [7 : 0] s_axi_awlen
          .s_axi_awsize(fsimtop_s_1_axi_awsize),      // input wire [2 : 0] s_axi_awsize
          .s_axi_awburst(fsimtop_s_1_axi_awburst),    // input wire [1 : 0] s_axi_awburst
          .s_axi_awlock(fsimtop_s_1_axi_awlock),      // input wire [0 : 0] s_axi_awlock
          // CACHE = xx1x indicates the transcation is modifiable and
          // that the converter should pack narrow writes into wider ones
          .s_axi_awcache(4'h2),    // input wire [3 : 0] s_axi_awcache
          .s_axi_awprot(fsimtop_s_1_axi_awprot),      // input wire [2 : 0] s_axi_awprot
          .s_axi_awregion(fsimtop_s_1_axi_awregion),  // input wire [3 : 0] s_axi_awregion
          .s_axi_awqos(fsimtop_s_1_axi_awqos),        // input wire [3 : 0] s_axi_awqos
          .s_axi_awvalid(fsimtop_s_1_axi_awvalid),    // input wire s_axi_awvalid
          .s_axi_awready(fsimtop_s_1_axi_awready),    // output wire s_axi_awready

          .s_axi_wdata(fsimtop_s_1_axi_wdata),        // input wire [63 : 0] s_axi_wdata
          .s_axi_wstrb(fsimtop_s_1_axi_wstrb),        // input wire [7 : 0] s_axi_wstrb
          .s_axi_wlast(fsimtop_s_1_axi_wlast),        // input wire s_axi_wlast
          .s_axi_wvalid(fsimtop_s_1_axi_wvalid),      // input wire s_axi_wvalid
          .s_axi_wready(fsimtop_s_1_axi_wready),      // output wire s_axi_wready

          .s_axi_bid(fsimtop_s_1_axi_bid),            // output wire [15 : 0] s_axi_bid
          .s_axi_bresp(fsimtop_s_1_axi_bresp),        // output wire [1 : 0] s_axi_bresp
          .s_axi_bvalid(fsimtop_s_1_axi_bvalid),      // output wire s_axi_bvalid
          .s_axi_bready(fsimtop_s_1_axi_bready),      // input wire s_axi_bready

          .s_axi_arid(fsimtop_s_1_axi_arid),          // input wire [15 : 0] s_axi_arid
          .s_axi_araddr(fsimtop_s_1_axi_araddr),      // input wire [63 : 0] s_axi_araddr
          .s_axi_arlen(fsimtop_s_1_axi_arlen),        // input wire [7 : 0] s_axi_arlen
          .s_axi_arsize(fsimtop_s_1_axi_arsize),      // input wire [2 : 0] s_axi_arsize
          .s_axi_arburst(fsimtop_s_1_axi_arburst),    // input wire [1 : 0] s_axi_arburst
          .s_axi_arlock(fsimtop_s_1_axi_arlock),      // input wire [0 : 0] s_axi_arlock
          // CACHE = xx1x indicates the transcation is modifiable and
          // that the converter should pack narrow reads into wider ones
          .s_axi_arcache(4'h2),                     // input wire [3 : 0] s_axi_arcache
          .s_axi_arprot(fsimtop_s_1_axi_arprot),      // input wire [2 : 0] s_axi_arprot
          .s_axi_arregion(fsimtop_s_1_axi_arregion),  // input wire [3 : 0] s_axi_arregion
          .s_axi_arqos(fsimtop_s_1_axi_arqos),        // input wire [3 : 0] s_axi_arqos
          .s_axi_arvalid(fsimtop_s_1_axi_arvalid),    // input wire s_axi_arvalid
          .s_axi_arready(fsimtop_s_1_axi_arready),    // output wire s_axi_arready

          .s_axi_rid(fsimtop_s_1_axi_rid),            // output wire [15 : 0] s_axi_rid
          .s_axi_rdata(fsimtop_s_1_axi_rdata),        // output wire [63 : 0] s_axi_rdata
          .s_axi_rresp(fsimtop_s_1_axi_rresp),        // output wire [1 : 0] s_axi_rresp
          .s_axi_rlast(fsimtop_s_1_axi_rlast),        // output wire s_axi_rlast
          .s_axi_rvalid(fsimtop_s_1_axi_rvalid),      // output wire s_axi_rvalid
          .s_axi_rready(fsimtop_s_1_axi_rready),      // input wire s_axi_rready

          .m_axi_aclk(clk),          // input wire m_axi_aclk
          .m_axi_aresetn(rst_main_n_sync),    // input wire m_axi_aresetn

          .m_axi_awid(clock_converted_axi_1_awid),          // output wire [15 : 0] m_axi_awid
          .m_axi_awaddr(clock_converted_axi_1_awaddr),      // output wire [63 : 0] m_axi_awaddr
          .m_axi_awlen(clock_converted_axi_1_awlen),        // output wire [7 : 0] m_axi_awlen
          .m_axi_awsize(clock_converted_axi_1_awsize),      // output wire [2 : 0] m_axi_awsize
          .m_axi_awburst(clock_converted_axi_1_awburst),    // output wire [1 : 0] m_axi_awburst
          .m_axi_awlock(clock_converted_axi_1_awlock),      // output wire [0 : 0] m_axi_awlock
          .m_axi_awcache(clock_converted_axi_1_awcache),    // output wire [3 : 0] m_axi_awcache
          .m_axi_awprot(clock_converted_axi_1_awprot),      // output wire [2 : 0] m_axi_awprot
          .m_axi_awregion(clock_converted_axi_1_awregion),  // output wire [3 : 0] m_axi_awregion
          .m_axi_awqos(clock_converted_axi_1_awqos),        // output wire [3 : 0] m_axi_awqos
          .m_axi_awvalid(clock_converted_axi_1_awvalid),    // output wire m_axi_awvalid
          .m_axi_awready(clock_converted_axi_1_awready),    // input wire m_axi_awready

          .m_axi_wdata(clock_converted_axi_1_wdata),        // output wire [511 : 0] m_axi_wdata
          .m_axi_wstrb(clock_converted_axi_1_wstrb),        // output wire [63 : 0] m_axi_wstrb
          .m_axi_wlast(clock_converted_axi_1_wlast),        // output wire m_axi_wlast
          .m_axi_wvalid(clock_converted_axi_1_wvalid),      // output wire m_axi_wvalid
          .m_axi_wready(clock_converted_axi_1_wready),      // input wire m_axi_wready

          .m_axi_bid(clock_converted_axi_1_bid),            // input wire [15 : 0] m_axi_bid
          .m_axi_bresp(clock_converted_axi_1_bresp),        // input wire [1 : 0] m_axi_bresp
          .m_axi_bvalid(clock_converted_axi_1_bvalid),      // input wire m_axi_bvalid
          .m_axi_bready(clock_converted_axi_1_bready),      // output wire m_axi_bready

          .m_axi_arid(clock_converted_axi_1_arid),          // output wire [15 : 0] m_axi_arid
          .m_axi_araddr(clock_converted_axi_1_araddr),      // output wire [63 : 0] m_axi_araddr
          .m_axi_arlen(clock_converted_axi_1_arlen),        // output wire [7 : 0] m_axi_arlen
          .m_axi_arsize(clock_converted_axi_1_arsize),      // output wire [2 : 0] m_axi_arsize
          .m_axi_arburst(clock_converted_axi_1_arburst),    // output wire [1 : 0] m_axi_arburst
          .m_axi_arlock(clock_converted_axi_1_arlock),      // output wire [0 : 0] m_axi_arlock
          .m_axi_arcache(clock_converted_axi_1_arcache),    // output wire [3 : 0] m_axi_arcache
          .m_axi_arprot(clock_converted_axi_1_arprot),      // output wire [2 : 0] m_axi_arprot
          .m_axi_arregion(clock_converted_axi_1_arregion),  // output wire [3 : 0] m_axi_arregion
          .m_axi_arqos(clock_converted_axi_1_arqos),        // output wire [3 : 0] m_axi_arqos
          .m_axi_arvalid(clock_converted_axi_1_arvalid),    // output wire m_axi_arvalid
          .m_axi_arready(clock_converted_axi_1_arready),    // input wire m_axi_arready

          .m_axi_rid(clock_converted_axi_1_rid),            // input wire [15 : 0] m_axi_rid
          .m_axi_rdata(clock_converted_axi_1_rdata),        // input wire [511 : 0] m_axi_rdata
          .m_axi_rresp(clock_converted_axi_1_rresp),        // input wire [1 : 0] m_axi_rresp
          .m_axi_rlast(clock_converted_axi_1_rlast),        // input wire m_axi_rlast
          .m_axi_rvalid(clock_converted_axi_1_rvalid),      // input wire m_axi_rvalid
          .m_axi_rready(clock_converted_axi_1_rready)      // output wire m_axi_rready
        );

        /* steps to move:
         * 1) copy clock converter's M interfaces to dwidth converter's M interfaces: DONE
         * 2) create clock_converted_* signals for clock M to width adapt S: DONE
         * 3) add asserts on arsize and awsize to confirm that they're always b110
        */

        assign DDRB_M_AXI_awid = 16'b0; // dwidth convert has no awid for some reason...
        assign DDRB_M_AXI_arid = 16'b0; // dwidth convert has no arid for some reason...
        // unused: DDRB_M_AXI_bid
        // unused: DDRB_M_AXI_rid

        axi_dwidth_converter_0 dwidth_adapt_64bits_512bits_1 (
          .s_axi_aclk(clk),          // input wire s_axi_aclk
          .s_axi_aresetn(rst_main_n_sync),    // input wire s_axi_aresetn

          .s_axi_awid(clock_converted_axi_1_awid),          // input wire [15 : 0] s_axi_awid
          .s_axi_awaddr(clock_converted_axi_1_awaddr),      // input wire [63 : 0] s_axi_awaddr
          .s_axi_awlen(clock_converted_axi_1_awlen),        // input wire [7 : 0] s_axi_awlen
          .s_axi_awsize(clock_converted_axi_1_awsize),      // input wire [2 : 0] s_axi_awsize
          .s_axi_awburst(clock_converted_axi_1_awburst),    // input wire [1 : 0] s_axi_awburst
          .s_axi_awlock(clock_converted_axi_1_awlock),      // input wire [0 : 0] s_axi_awlock
          .s_axi_awcache(clock_converted_axi_1_awcache),    // input wire [3 : 0] s_axi_awcache
          .s_axi_awprot(clock_converted_axi_1_awprot),      // input wire [2 : 0] s_axi_awprot
          .s_axi_awregion(clock_converted_axi_1_awregion),  // input wire [3 : 0] s_axi_awregion
          .s_axi_awqos(clock_converted_axi_1_awqos),        // input wire [3 : 0] s_axi_awqos
          .s_axi_awvalid(clock_converted_axi_1_awvalid),    // input wire s_axi_awvalid
          .s_axi_awready(clock_converted_axi_1_awready),    // output wire s_axi_awready

          .s_axi_wdata(clock_converted_axi_1_wdata),        // input wire [63 : 0] s_axi_wdata
          .s_axi_wstrb(clock_converted_axi_1_wstrb),        // input wire [7 : 0] s_axi_wstrb
          .s_axi_wlast(clock_converted_axi_1_wlast),        // input wire s_axi_wlast
          .s_axi_wvalid(clock_converted_axi_1_wvalid),      // input wire s_axi_wvalid
          .s_axi_wready(clock_converted_axi_1_wready),      // output wire s_axi_wready

          .s_axi_bid(clock_converted_axi_1_bid),            // output wire [15 : 0] s_axi_bid
          .s_axi_bresp(clock_converted_axi_1_bresp),        // output wire [1 : 0] s_axi_bresp
          .s_axi_bvalid(clock_converted_axi_1_bvalid),      // output wire s_axi_bvalid
          .s_axi_bready(clock_converted_axi_1_bready),      // input wire s_axi_bready

          .s_axi_arid(clock_converted_axi_1_arid),          // input wire [15 : 0] s_axi_arid
          .s_axi_araddr(clock_converted_axi_1_araddr),      // input wire [63 : 0] s_axi_araddr
          .s_axi_arlen(clock_converted_axi_1_arlen),        // input wire [7 : 0] s_axi_arlen
          .s_axi_arsize(clock_converted_axi_1_arsize),      // input wire [2 : 0] s_axi_arsize
          .s_axi_arburst(clock_converted_axi_1_arburst),    // input wire [1 : 0] s_axi_arburst
          .s_axi_arlock(clock_converted_axi_1_arlock),      // input wire [0 : 0] s_axi_arlock
          .s_axi_arcache(clock_converted_axi_1_arcache),    // input wire [3 : 0] s_axi_arcache
          .s_axi_arprot(clock_converted_axi_1_arprot),      // input wire [2 : 0] s_axi_arprot
          .s_axi_arregion(clock_converted_axi_1_arregion),  // input wire [3 : 0] s_axi_arregion
          .s_axi_arqos(clock_converted_axi_1_arqos),        // input wire [3 : 0] s_axi_arqos
          .s_axi_arvalid(clock_converted_axi_1_arvalid),    // input wire s_axi_arvalid
          .s_axi_arready(clock_converted_axi_1_arready),    // output wire s_axi_arready

          .s_axi_rid(clock_converted_axi_1_rid),            // output wire [15 : 0] s_axi_rid
          .s_axi_rdata(clock_converted_axi_1_rdata),        // output wire [63 : 0] s_axi_rdata
          .s_axi_rresp(clock_converted_axi_1_rresp),        // output wire [1 : 0] s_axi_rresp
          .s_axi_rlast(clock_converted_axi_1_rlast),        // output wire s_axi_rlast
          .s_axi_rvalid(clock_converted_axi_1_rvalid),      // output wire s_axi_rvalid
          .s_axi_rready(clock_converted_axi_1_rready),      // input wire s_axi_rready


          .m_axi_awaddr(DDRB_M_AXI_awaddr),      // output wire [63 : 0] m_axi_awaddr
          .m_axi_awlen(DDRB_M_AXI_awlen),        // output wire [7 : 0] m_axi_awlen
          .m_axi_awsize(DDRB_M_AXI_awsize),      // output wire [2 : 0] m_axi_awsize
          .m_axi_awburst(DDRB_M_AXI_awburst),    // output wire [1 : 0] m_axi_awburst
          .m_axi_awlock(DDRB_M_AXI_awlock),      // output wire [0 : 0] m_axi_awlock
          .m_axi_awcache(DDRB_M_AXI_awcache),    // output wire [3 : 0] m_axi_awcache
          .m_axi_awprot(DDRB_M_AXI_awprot),      // output wire [2 : 0] m_axi_awprot
          .m_axi_awregion(DDRB_M_AXI_awregion),  // output wire [3 : 0] m_axi_awregion
          .m_axi_awqos(DDRB_M_AXI_awqos),        // output wire [3 : 0] m_axi_awqos
          .m_axi_awvalid(DDRB_M_AXI_awvalid),    // output wire m_axi_awvalid
          .m_axi_awready(DDRB_M_AXI_awready),    // input wire m_axi_awready

          .m_axi_wdata(DDRB_M_AXI_wdata),        // output wire [511 : 0] m_axi_wdata
          .m_axi_wstrb(DDRB_M_AXI_wstrb),        // output wire [63 : 0] m_axi_wstrb
          .m_axi_wlast(DDRB_M_AXI_wlast),        // output wire m_axi_wlast
          .m_axi_wvalid(DDRB_M_AXI_wvalid),      // output wire m_axi_wvalid
          .m_axi_wready(DDRB_M_AXI_wready),      // input wire m_axi_wready

          .m_axi_bresp(DDRB_M_AXI_bresp),        // input wire [1 : 0] m_axi_bresp
          .m_axi_bvalid(DDRB_M_AXI_bvalid),      // input wire m_axi_bvalid
          .m_axi_bready(DDRB_M_AXI_bready),      // output wire m_axi_bready

          .m_axi_araddr(DDRB_M_AXI_araddr),      // output wire [63 : 0] m_axi_araddr
          .m_axi_arlen(DDRB_M_AXI_arlen),        // output wire [7 : 0] m_axi_arlen
          .m_axi_arsize(DDRB_M_AXI_arsize),      // output wire [2 : 0] m_axi_arsize
          .m_axi_arburst(DDRB_M_AXI_arburst),    // output wire [1 : 0] m_axi_arburst
          .m_axi_arlock(DDRB_M_AXI_arlock),      // output wire [0 : 0] m_axi_arlock
          .m_axi_arcache(DDRB_M_AXI_arcache),    // output wire [3 : 0] m_axi_arcache
          .m_axi_arprot(DDRB_M_AXI_arprot),      // output wire [2 : 0] m_axi_arprot
          .m_axi_arregion(DDRB_M_AXI_arregion),  // output wire [3 : 0] m_axi_arregion
          .m_axi_arqos(DDRB_M_AXI_arqos),        // output wire [3 : 0] m_axi_arqos
          .m_axi_arvalid(DDRB_M_AXI_arvalid),    // output wire m_axi_arvalid
          .m_axi_arready(DDRB_M_AXI_arready),    // input wire m_axi_arready

          .m_axi_rdata(DDRB_M_AXI_rdata),        // input wire [511 : 0] m_axi_rdata
          .m_axi_rresp(DDRB_M_AXI_rresp),        // input wire [1 : 0] m_axi_rresp
          .m_axi_rlast(DDRB_M_AXI_rlast),        // input wire m_axi_rlast
          .m_axi_rvalid(DDRB_M_AXI_rvalid),      // input wire m_axi_rvalid
          .m_axi_rready(DDRB_M_AXI_rready)      // output wire m_axi_rready
        );
    end
    else begin
        assign DDRB_M_AXI_awaddr = '0;
        assign DDRB_M_AXI_awlen = '0;
        assign DDRB_M_AXI_awsize = '0;
        assign DDRB_M_AXI_awburst = '0;
        assign DDRB_M_AXI_awid = '0;
        assign DDRB_M_AXI_awvalid = '0;
        assign DDRB_M_AXI_awready = '0;

        assign DDRB_M_AXI_wdata = '0;
        assign DDRB_M_AXI_wstrb = '0;
        assign DDRB_M_AXI_wlast = '0;
        assign DDRB_M_AXI_wvalid = '0;
        assign DDRB_M_AXI_wready = '0;

        assign DDRB_M_AXI_bready = '0;

        assign DDRB_M_AXI_arid = '0;
        assign DDRB_M_AXI_araddr = '0;
        assign DDRB_M_AXI_arlen = '0;
        assign DDRB_M_AXI_arsize = '0;
        assign DDRB_M_AXI_arburst = '0;
        assign DDRB_M_AXI_arvalid = '0;

        assign DDRB_M_AXI_rready = '0;


        assign fsimtop_s_1_axi_awready = '0;
        assign fsimtop_s_1_axi_wready = '0;
        assign fsimtop_s_1_axi_arready = '0;

        assign fsimtop_s_1_axi_bid = '0;
        assign fsimtop_s_1_axi_bresp = '0;
        assign fsimtop_s_1_axi_bvalid = '0;

        assign fsimtop_s_1_axi_rid = '0;
        assign fsimtop_s_1_axi_rdata = '0;
        assign fsimtop_s_1_axi_rresp = '0;
        assign fsimtop_s_1_axi_rlast = '0;
        assign fsimtop_s_1_axi_rvalid = '0;
    end
endgenerate

endmodule
